module xor_gate (input i_a, input i_b, output o_f);

   assign o_f = i_a ^ i_b;

endmodule
