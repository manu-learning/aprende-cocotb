module xor_gate (input entrada_A, input entrada_B, output salida_F);

   assign salida_F = entrada_A ^ entrada_B;

endmodule
